----------------------------------------------------------------------------------
-- Sourced from: vhdlguru, pwkolas
-- URL: https://vhdlguru.blogspot.com/2017/09/pushbutton-debounce-circuit-in-vhdl.html
-- Modified by: Jeremy, Randipa, Geeth
-- Create Date: 13.05.2020 22:14:45
-- Design Name: 
-- Module Name: button_debouncer - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity btn_debouncer is
    port(   Clock : in std_logic;
            Reset : in std_logic := '0';
            button_in : in std_logic;
            pulse_out : out std_logic
        );
end btn_debouncer;

architecture behav of btn_debouncer is

--the below constants decide the working parameters.
--the higher this is, the more longer time the user has to press the button.
constant COUNT_MAX : integer := 250; 
--set it '1' if the button creates a high pulse when its pressed, otherwise '0'.
constant BTN_ACTIVE : std_logic := '1';

signal count : integer := 0;
type state_type is (idle,wait_time); --state machine
signal state : state_type := idle;

begin
  
process(Reset,Clock)
begin
    --Asynchronous reset
    if(Reset = '1') then
        state <= idle;
        pulse_out <= '0';
   --Counting up in the rising edge
   elsif(rising_edge(Clock)) then
        case (state) is
            when idle =>
                if(button_in = BTN_ACTIVE) then  
                    state <= wait_time;
                else
                    state <= idle; --wait until button is pressed.
                end if;
                pulse_out <= '0';
            when wait_time =>
                if(count = COUNT_MAX) then
                    count <= 0;
                    if(button_in = BTN_ACTIVE) then
                        pulse_out <= '1';
                    end if;
                    state <= idle;  
                else
                    count <= count + 1;
                end if; 
        end case;       
    end if;        
end process;                  
                                                                                
end architecture behav;